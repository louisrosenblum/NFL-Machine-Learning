A.J. Brown,25.4,22,15,10,76,48,927,19.3,7,36,91,3.2,61.8,63.20%,12.2,3,60,1,2,49,20,4,0.2,51,19.4,987,0.40,0.07,0.17,0.00,20.67,12.27,166.47,13.57,1.13,0.00
Aaron Jones,17.1,25,15,15,62,47,431,9.2,3,16,67,3.1,28.7,75.80%,7,211,984,16,50,56,4.7,65.6,14.1,258,5.5,1415,23.07,84.67,3.67,0.93,7.20,5.47,38.40,7.02,0.13,0.07
Adam Thielen,6,29,10,10,48,30,418,13.9,6,18,44,3,41.8,62.50%,8.7,4,6,1,1,3,1.5,0.6,0.4,34,12.5,424,0.53,2.00,3.75,0.00,15.47,11.07,129.33,11.69,0.67,0.00
Adrian Peterson,18.1,34,14,14,19,16,142,8.9,0,7,22,1.1,10.1,84.20%,7.5,198,820,5,38,29,4.1,58.6,14.1,214,4.5,962,18.73,67.80,3.62,0.60,7.47,5.53,40.73,7.36,0.07,0.13
Albert Wilson,10.9,27,12,3,54,38,292,7.7,1,18,35,3.2,24.3,70.40%,5.4,5,45,0,1,28,9,3.8,0.4,43,7.8,337,0.33,1.73,5.20,0.00,19.60,13.13,186.47,14.20,1.47,0.13
Alec Ingold,5.2,23,15,4,6,6,44,7.3,1,4,14,0.4,2.9,100.00%,7.3,9,17,0,7,4,1.9,1.1,0.6,15,4.1,61,22.33,119.13,5.33,1.07,6.60,5.33,49.87,9.35,0.27,0.13
Alex Armah,0,25,15,1,2,2,6,3,0,0,4,0.1,0.4,100.00%,3,6,11,1,1,4,1.8,0.7,0.4,8,2.1,17,19.27,82.27,4.27,1.07,6.80,5.53,49.67,8.98,0.07,0.33
Alex Erickson,-0.4,27,15,5,74,42,513,12.2,0,25,52,2.8,34.2,56.80%,6.9,4,28,0,2,17,7,1.9,0.3,46,11.8,541,0.33,4.80,14.40,0.07,19.87,9.93,117.60,11.84,0.27,0.20
Alfred Morris,0,31,1,0,0,0,0,,0,0,0,0,0,0.00%,,1,4,0,1,4,4,4,1,1,4,4,21.80,106.53,4.89,0.80,5.87,4.67,42.87,9.19,0.27,0.20
Allen Hurns,1.9,28,14,7,47,32,416,13,2,18,27,2.3,29.7,68.10%,8.9,,,,0,,,,,32,13,416,0.33,1.73,5.20,0.00,19.60,13.13,186.47,14.20,1.47,0.13
Allen Lazard,3.4,24,15,2,44,31,408,13.2,2,20,43,2.1,27.2,70.50%,9.3,1,21,0,1,21,21,1.4,0.1,32,13.4,429,0.20,1.13,5.67,0.00,18.93,11.47,147.87,12.90,0.60,0.13
Allen Robinson,19.5,26,15,14,142,89,1076,12.1,7,57,49,5.9,71.7,62.70%,7.6,,,,0,,,,,89,12.1,1076,0.47,1.40,3.00,0.00,17.67,10.00,159.13,15.91,0.73,0.07
Alvin Kamara,13.9,24,13,9,94,79,515,6.5,1,27,41,6.1,39.6,84.00%,5.5,163,758,3,29,40,4.7,58.3,12.5,242,5.3,1273,20.13,83.87,4.17,0.27,7.80,6.73,45.33,6.73,0.13,0.27
Amari Cooper,2.9,25,15,15,114,75,1097,14.6,8,51,53,5,73.1,65.80%,9.6,,,,0,,,,,75,14.6,1097,0.53,1.80,3.38,0.07,19.93,12.53,151.60,12.10,0.80,0.27
Ameer Abdullah,2.5,26,15,0,17,12,74,6.2,1,5,16,0.8,4.9,70.60%,4.4,17,93,0,3,15,5.5,6.2,1.1,29,5.8,167,23.07,94.20,4.08,0.80,7.07,5.60,40.07,7.15,0.27,0.00
Andre Patton,1.8,25,12,4,14,6,56,9.3,0,4,15,0.5,4.7,42.90%,4,,,,0,,,,,6,9.3,56,0.60,2.00,3.33,0.00,21.27,14.33,171.60,11.97,1.20,0.27
Andre Roberts,1.7,31,13,0,7,3,20,6.7,0,1,7,0.2,1.5,42.90%,2.9,1,7,0,0,7,7,0.5,0.1,4,6.8,27,0.33,2.60,7.80,0.00,18.80,11.07,145.73,13.17,0.87,0.20
Andrew Beck,3.3,23,15,5,10,7,82,11.7,0,5,29,0.5,5.5,70.00%,8.2,1,3,0,1,3,3,0.2,0.1,8,10.6,85,22.20,108.87,4.90,0.60,8.00,5.67,55.47,9.79,0.33,0.20
Andy Isabella,1.3,23,14,1,13,9,189,21,1,4,88,0.6,13.5,69.20%,14.5,4,15,0,0,6,3.8,1.1,0.3,13,15.7,204,0.87,7.13,8.23,0.00,18.47,11.27,144.00,12.78,0.73,0.07
Anthony Firkser,1.7,24,14,1,22,13,199,15.3,1,9,39,0.9,14.2,59.10%,9,,,,0,,,,,13,15.3,199,0.07,3.80,57.00,0.00,7.47,4.87,58.60,12.04,0.33,0.00
Anthony Miller,26.8,25,15,6,84,51,651,12.8,2,34,35,3.4,43.4,60.70%,7.8,1,-1,0,0,-1,-1,-0.1,0.1,52,12.5,650,0.47,1.40,3.00,0.00,17.67,10.00,159.13,15.91,0.73,0.07
Anthony Sherman,0,31,15,0,3,2,22,11,0,2,15,0.1,1.5,66.70%,7.3,4,9,0,3,5,2.3,0.6,0.3,6,5.2,31,23.73,94.00,3.96,0.47,6.53,5.20,34.80,6.69,0.13,0.20
Antonio Callaway,0,22,4,2,15,8,89,11.1,0,3,41,2,22.3,53.30%,5.9,,,,0,,,,,8,11.1,89,0.33,2.80,8.40,0.00,20.33,13.87,170.33,12.28,0.93,0.07
Ashton Dulin,1.4,22,12,0,2,2,17,8.5,0,0,13,0.2,1.4,100.00%,8.5,,,,0,,,,,2,8.5,17,1.27,13.80,10.89,0.07,21.20,12.67,175.80,13.88,1.20,0.13
Austin Ekeler,13.1,24,15,8,97,83,950,11.4,8,40,84,5.5,63.3,85.60%,9.8,123,511,3,29,35,4.2,34.1,8.2,206,7.1,1461,22.13,96.27,4.35,0.47,6.53,4.67,36.13,7.74,0.27,0.27
Austin Hooper,5,25,12,9,88,68,742,10.9,6,38,35,5.7,61.8,77.30%,8.4,,,,0,,,,,68,10.9,742,0.00,0.00,0.00,0.00,6.07,4.07,34.80,8.56,0.40,0.07
Ben Koyack,0,26,10,5,3,1,9,9,0,0,9,0.1,0.9,33.30%,3,,,,0,,,,,1,9,9,0.07,-0.33,-5.00,0.00,7.20,4.60,57.07,12.41,0.60,0.00
Ben Watson,0,39,9,7,23,16,169,10.6,0,9,26,1.8,18.8,69.60%,7.3,,,,0,,,,,16,10.6,169,0.13,0.47,3.50,0.00,6.27,4.40,53.20,12.09,0.40,0.07
Bennie Fowler,0,28,8,2,36,23,193,8.4,0,12,17,2.9,24.1,63.90%,5.4,1,20,0,1,20,20,2.5,0.1,24,8.9,213,0.53,1.80,3.38,0.00,20.80,12.33,179.00,14.51,1.80,0.00
Benny Snell,0.1,21,12,1,4,3,23,7.7,0,0,14,0.3,1.9,75.00%,5.8,90,335,1,15,23,3.7,27.9,7.5,93,3.8,358,19.93,89.27,4.48,0.60,7.47,5.47,42.33,7.74,0.20,0.13
Blake Bell,6.1,28,14,7,13,7,66,9.4,0,3,30,0.5,4.7,53.80%,5.1,,,,0,,,,,7,9.4,66,0.00,0.00,0.00,0.00,7.87,5.53,57.53,10.40,0.20,0.00
Blake Jarwin,6,25,15,7,40,31,365,11.8,3,17,42,2.1,24.3,77.50%,9.1,,,,0,,,,,31,11.8,365,0.13,0.60,4.50,0.00,6.53,4.33,52.93,12.22,0.33,0.00
Bobo Wilson,0,24,6,1,11,3,35,11.7,0,2,14,0.5,5.8,27.30%,3.2,,,,0,,,,,3,11.7,35,0.33,1.73,5.20,0.00,22.47,13.73,188.73,13.74,1.20,0.27
Boston Scott,13.5,24,10,2,20,20,120,6,0,7,17,2,12,100.00%,6,42,191,2,12,25,4.5,19.1,4.2,62,5,311,25.80,119.33,4.63,0.67,7.73,6.07,53.13,8.76,0.27,0.20
Brandin Cooks,8.6,26,13,13,67,39,543,13.9,2,29,57,3,41.8,58.20%,8.1,6,52,0,3,27,8.7,4,0.5,45,13.2,595,0.67,3.27,4.90,0.00,17.67,10.87,135.47,12.47,0.80,0.00
Brandon Bolden,0,29,14,2,11,9,111,12.3,1,6,29,0.6,7.9,81.80%,10.1,15,68,3,5,21,4.5,4.9,1.1,24,7.5,179,24.87,115.73,4.65,0.80,5.87,4.80,44.20,9.21,0.27,0.20
Brandon Zylstra,0,26,7,0,4,2,10,5,0,1,7,0.3,1.4,50.00%,2.5,,,,0,,,,,2,5,10,1.27,11.87,9.37,0.00,21.53,12.73,157.27,12.35,0.80,0.13
Braxton Berrios,0,24,15,0,11,5,104,20.8,0,2,69,0.3,6.9,45.50%,9.5,,,,0,,,,,5,20.8,104,0.47,3.73,8.00,0.00,22.60,13.33,166.27,12.47,0.73,0.27
Breshad Perriman,34.6,26,13,3,61,31,511,16.5,5,24,44,2.4,39.3,50.80%,8.4,2,16,0,1,13,8,1.2,0.2,33,16,527,0.33,1.73,5.20,0.00,22.47,13.73,188.73,13.74,1.20,0.27
Brian Hill,1.6,24,11,2,14,10,69,6.9,1,4,12,0.9,6.3,71.40%,4.9,73,302,2,18,27,4.1,27.5,6.6,83,4.5,371,19.27,80.87,4.20,0.40,5.53,3.87,24.67,6.38,0.00,0.33
Buddy Howell,0,23,15,0,0,0,0,,0,0,0,0,0,0.00%,,2,5,0,0,4,2.5,0.3,0.1,2,2.5,5,21.60,87.07,4.03,0.80,8.20,6.33,46.87,7.40,0.20,0.13
Byron Pringle,0,26,15,0,16,12,170,14.2,1,7,28,0.8,11.3,75.00%,10.6,,,,0,,,,,12,14.2,170,0.53,5.93,11.12,0.00,17.00,10.53,136.40,12.95,0.87,0.07
C.J. Anderson,0,28,2,0,0,0,0,,0,0,0,0,0,0.00%,,16,43,0,1,9,2.7,21.5,8,16,2.7,43,18.13,54.67,3.01,0.53,7.27,5.40,31.00,5.74,0.07,0.40
C.J. Board,1.8,26,3,0,4,2,31,15.5,0,1,23,0.7,10.3,50.00%,7.8,,,,0,,,,,2,15.5,31,0.67,4.07,6.10,0.07,17.67,10.93,170.00,15.55,1.13,0.07
C.J. Ham,4.8,26,15,7,25,17,149,8.8,1,6,36,1.1,9.9,68.00%,6,5,13,0,1,9,2.6,0.9,0.3,22,7.4,162,23.07,94.20,4.08,0.80,7.07,5.60,40.07,7.15,0.27,0.00
C.J. Prosise,3.5,25,9,0,12,10,76,7.6,0,3,21,1.1,8.4,83.30%,6.3,23,72,1,4,17,3.1,8,2.6,33,4.5,148,23.40,127.27,5.44,1.67,5.07,3.80,23.47,6.18,0.20,0.07
C.J. Uzomah,1.8,26,15,15,34,22,217,9.9,1,10,36,1.5,14.5,64.70%,6.4,,,,0,,,,,22,9.9,217,0.07,0.27,4.00,0.07,5.80,3.80,42.20,11.11,0.27,0.07
Cameron Brate,6.3,28,15,6,52,35,309,8.8,3,20,37,2.3,20.6,67.30%,5.9,,,,0,,,,,35,8.8,309,0.13,2.00,15.00,0.00,6.47,4.60,51.53,11.20,0.33,0.00
Carlos Hyde,16.4,29,15,13,16,10,42,4.2,0,2,14,0.7,2.8,62.50%,2.6,241,1057,6,54,58,4.4,70.5,16.1,251,4.4,1099,21.60,87.07,4.03,0.80,8.20,6.33,46.87,7.40,0.20,0.13
Charles Clay,2.8,30,15,10,24,18,237,13.2,1,12,47,1.2,15.8,75.00%,9.9,,,,0,,,,,18,13.2,237,0.13,1.87,14.00,0.00,6.33,4.20,49.80,11.86,0.60,0.00
Chase Edmonds,0,23,12,2,21,12,105,8.8,1,5,31,1,8.8,57.10%,5,59,304,4,12,37,5.2,25.3,4.9,71,5.8,409,21.80,106.53,4.89,0.80,5.87,4.67,42.87,9.19,0.27,0.20
Chris Carson,26.7,25,15,15,47,37,266,7.2,2,10,21,2.5,17.7,78.70%,5.7,278,1230,7,75,59,4.4,82,18.5,315,4.7,1496,23.40,127.27,5.44,1.67,5.07,3.80,23.47,6.18,0.20,0.07
Chris Conley,20.9,27,15,13,84,44,737,16.8,5,34,70,2.9,49.1,52.40%,8.8,,,,0,,,,,44,16.8,737,0.67,4.07,6.10,0.07,17.67,10.93,170.00,15.55,1.13,0.07
Chris Hogan,2.3,32,6,0,11,6,53,8.8,0,2,13,1,8.8,54.50%,4.8,,,,0,,,,,6,8.8,53,1.27,11.87,9.37,0.00,21.53,12.73,157.27,12.35,0.80,0.13
Chris Manhertz,0,27,14,5,1,1,11,11,0,1,11,0.1,0.8,100.00%,11,,,,0,,,,,1,11,11,0.00,0.00,0.00,0.00,8.73,6.00,67.53,11.26,0.40,0.07
Chris Moore,0,26,13,1,5,3,21,7,0,0,13,0.2,1.6,60.00%,4.2,,,,0,,,,,3,7,21,0.47,2.20,4.71,0.00,20.87,13.13,164.20,12.50,1.33,0.13
Chris Thompson,4.6,29,10,0,55,41,378,9.2,0,16,39,4.1,37.8,74.50%,6.9,34,127,0,6,12,3.7,12.7,3.4,75,6.7,505,18.73,67.80,3.62,0.60,7.47,5.53,40.73,7.36,0.07,0.13
Christian Blake,0,23,8,2,22,11,91,8.3,0,5,13,1.4,11.4,50.00%,4.1,,,,0,,,,,11,8.3,91,1.13,7.53,6.65,0.07,19.27,11.53,129.13,11.20,1.00,0.27
Christian Kirk,10.1,23,12,12,98,61,649,10.6,3,29,69,5.1,54.1,62.20%,6.6,9,87,0,4,28,9.7,7.3,0.8,70,10.5,736,0.87,7.13,8.23,0.00,18.47,11.27,144.00,12.78,0.73,0.07
Clive Walford,5.4,28,7,3,8,4,57,14.3,0,4,19,0.6,8.1,50.00%,7.1,0,4,0,0,4,,0.6,0,4,15.3,61,0.07,0.13,2.00,0.00,6.80,4.40,47.33,10.76,0.47,0.00
Cody Core,0,25,15,0,5,3,28,9.3,0,2,11,0.2,1.9,60.00%,5.6,,,,0,,,,,3,9.3,28,0.53,1.80,3.38,0.00,20.80,12.33,179.00,14.51,1.80,0.00
Cody Hollister,0,26,5,0,2,2,13,6.5,0,0,11,0.4,2.6,100.00%,6.5,,,,0,,,,,2,6.5,13,0.40,0.07,0.17,0.00,20.67,12.27,166.47,13.57,1.13,0.00
Cody Latimer,3.1,27,14,9,39,22,288,13.1,2,18,43,1.6,20.6,56.40%,7.4,,,,0,,,,,22,13.1,288,0.53,1.80,3.38,0.00,20.80,12.33,179.00,14.51,1.80,0.00
Cole Beasley,1.6,30,15,10,106,67,778,11.6,6,37,51,4.5,51.9,63.20%,7.3,,,,0,,,,,67,11.6,778,0.33,2.60,7.80,0.00,18.80,11.07,145.73,13.17,0.87,0.20
Cooper Kupp,16.1,26,15,13,124,87,1062,12.2,9,45,66,5.8,70.8,70.20%,8.6,2,4,0,0,6,2,0.3,0.1,89,12,1066,0.67,3.27,4.90,0.00,17.67,10.87,135.47,12.47,0.80,0.00
Corey Davis,8.7,24,14,10,64,39,557,14.3,2,29,38,2.8,39.8,60.90%,8.7,,,,0,,,,,39,14.3,557,0.40,0.07,0.17,0.00,20.67,12.27,166.47,13.57,1.13,0.00
Courtland Sutton,11.9,24,15,13,116,68,1060,15.6,6,47,70,4.5,70.7,58.60%,9.1,3,17,0,1,9,5.7,1.1,0.2,71,15.2,1077,0.40,3.33,8.33,0.00,17.20,9.53,122.40,12.84,0.67,0.07
Curtis Samuel,16.4,23,15,14,101,52,614,11.8,6,35,44,3.5,40.9,51.50%,6.1,19,130,1,7,16,6.8,8.7,1.3,71,10.5,744,1.27,11.87,9.37,0.00,21.53,12.73,157.27,12.35,0.80,0.13
D.J. Moore,20.3,22,15,15,135,87,1175,13.5,4,63,52,5.8,78.3,64.40%,8.7,6,40,0,3,13,6.7,2.7,0.4,93,13.1,1215,1.27,11.87,9.37,0.00,21.53,12.73,157.27,12.35,0.80,0.13
D.K. Metcalf,11.6,22,15,14,88,52,819,15.8,6,33,54,3.5,54.6,59.10%,9.3,2,11,0,0,7,5.5,0.7,0.1,54,15.4,830,0.40,3.40,8.50,0.07,22.20,14.47,180.60,12.48,0.80,0.07
DaeSean Hamilton,3.3,24,15,2,46,23,232,10.1,1,14,28,1.5,15.5,50.00%,5,,,,0,,,,,23,10.1,232,0.40,3.33,8.33,0.00,17.20,9.53,122.40,12.84,0.67,0.07
Dallas Goedert,10.5,24,14,8,77,54,542,10,5,30,28,3.9,38.7,70.10%,7,,,,0,,,,,54,10,542,0.13,0.00,0.00,0.00,7.67,5.47,57.27,10.48,0.60,0.00
Dalton Schultz,0,23,15,0,2,1,6,6,0,0,6,0.1,0.4,50.00%,3,,,,0,,,,,1,6,6,0.13,0.60,4.50,0.00,6.53,4.33,52.93,12.22,0.33,0.00
Dalyn Dawkins,0,25,2,0,1,0,0,,0,0,0,0,0,0.00%,0,11,26,0,2,14,2.4,13,5.5,11,2.4,26,20.67,90.87,4.40,0.40,8.07,6.87,58.93,8.58,0.53,0.07
Damiere Byrd,14.6,26,10,3,38,25,285,11.4,0,12,58,2.5,28.5,65.80%,7.5,,,,0,,,,,25,11.4,285,0.87,7.13,8.23,0.00,18.47,11.27,144.00,12.78,0.73,0.07
Damion Ratley,5.3,24,12,3,21,10,136,13.6,0,9,29,0.8,11.3,47.60%,6.5,,,,0,,,,,10,13.6,136,0.33,2.80,8.40,0.00,20.33,13.87,170.33,12.28,0.93,0.07
Dan Arnold,7.6,24,4,0,8,4,51,12.8,1,3,20,1,12.8,50.00%,6.4,,,,0,,,,,4,12.8,51,0.13,1.87,14.00,0.00,6.33,4.20,49.80,11.86,0.60,0.00
Daniel Brown,1.4,27,15,4,7,4,40,10,1,3,20,0.3,2.7,57.10%,5.7,,,,0,,,,,4,10,40,0.07,-0.20,-3.00,0.00,5.27,3.33,37.07,11.12,0.20,0.00
Danny Amendola,18.2,34,14,9,93,60,662,11,1,36,47,4.3,47.3,64.50%,7.1,,,,0,,,,,60,11,662,0.60,4.33,7.22,0.07,24.67,14.73,197.87,13.43,1.40,0.13
Danny Vitale,0,26,15,4,12,7,97,13.9,0,3,27,0.5,6.5,58.30%,8.1,1,3,0,0,3,3,0.2,0.1,8,12.5,100,23.07,84.67,3.67,0.93,7.20,5.47,38.40,7.02,0.13,0.07
Dante Pettis,0,24,11,4,24,11,109,9.9,2,7,21,1,9.9,45.80%,4.5,,,,0,,,,,11,9.9,109,0.73,2.93,4.00,0.00,17.60,11.93,164.93,13.82,1.00,0.20
Dare Ogunbowale,2.6,25,15,0,46,35,286,8.2,0,14,21,2.3,19.1,76.10%,6.2,10,13,2,3,12,1.3,0.9,0.7,45,6.6,299,24.33,98.53,4.05,0.87,6.93,5.20,54.40,10.46,0.53,0.33
Darius Jennings,0,27,7,0,5,2,17,8.5,0,2,11,0.3,2.4,40.00%,3.4,,,,0,,,,,2,8.5,17,0.40,0.07,0.17,0.00,20.67,12.27,166.47,13.57,1.13,0.00
Darius Slayton,11.1,22,13,9,75,44,690,15.7,8,31,55,3.4,53.1,58.70%,9.2,,,,0,,,,,44,15.7,690,0.53,1.80,3.38,0.00,20.80,12.33,179.00,14.51,1.80,0.00
Darrell Henderson,0,22,13,0,6,4,37,9.3,0,1,14,0.3,2.8,66.70%,6.2,39,147,0,10,22,3.8,11.3,3,43,4.3,184,20.40,81.40,3.99,0.73,7.93,6.13,47.00,7.66,0.13,0.13
Darren Fells,1.2,33,15,14,48,34,341,10,7,22,24,2.3,22.7,70.80%,7.1,,,,0,,,,,34,10,341,0.00,0.00,0.00,0.00,7.27,4.93,56.93,11.54,0.60,0.13
Darren Waller,20.2,27,15,15,107,84,1038,12.4,3,50,48,5.6,69.2,78.50%,9.7,2,5,0,0,7,2.5,0.3,0.1,86,12.1,1043,0.07,0.27,4.00,0.00,6.00,4.20,51.20,12.19,0.47,0.00
Darrius Shepherd,0,24,6,0,2,1,1,1,0,0,1,0.2,0.2,50.00%,0.5,,,,0,,,,,1,1,1,0.20,1.13,5.67,0.00,18.93,11.47,147.87,12.90,0.60,0.13
Darwin Thompson,4.9,23,11,0,9,8,47,5.9,0,2,19,0.7,4.3,88.90%,5.2,33,111,1,7,12,3.4,10.1,3,41,3.9,158,23.73,94.00,3.96,0.47,6.53,5.20,34.80,6.69,0.13,0.20
Davante Adams,23.3,27,11,11,114,76,904,11.9,4,49,58,6.9,82.2,66.70%,7.9,,,,0,,,,,76,11.9,904,0.20,1.13,5.67,0.00,18.93,11.47,147.87,12.90,0.60,0.13
David Johnson,0.6,28,13,9,47,36,370,10.3,4,17,31,2.8,28.5,76.60%,7.9,94,345,2,20,18,3.7,26.5,7.2,130,5.5,715,21.80,106.53,4.89,0.80,5.87,4.67,42.87,9.19,0.27,0.20
David Montgomery,5.9,22,15,8,35,25,185,7.4,1,7,30,1.7,12.3,71.40%,5.3,219,776,5,43,55,3.5,51.7,14.6,244,3.9,961,22.47,105.87,4.71,0.93,8.07,5.93,42.87,7.22,0.07,0.07
David Moore,0,24,13,1,32,15,271,18.1,2,12,60,1.2,20.8,46.90%,8.5,3,25,0,1,19,8.3,1.9,0.2,18,16.4,296,0.40,3.40,8.50,0.07,22.20,14.47,180.60,12.48,0.80,0.07
Dawson Knox,2.1,23,15,11,50,28,388,13.9,2,15,49,1.9,25.9,56.00%,7.8,1,9,0,1,9,9,0.6,0.1,29,13.7,397,0.00,0.00,0.00,0.00,5.93,4.13,41.87,10.13,0.53,0.00
DeAndre Carter,0,26,15,2,7,5,97,19.4,0,3,46,0.3,6.5,71.40%,13.9,,,,0,,,,,5,19.4,97,0.60,2.67,4.44,0.00,19.60,12.87,166.93,12.97,0.80,0.07
DeAndre Washington,4.2,26,15,2,32,28,237,8.5,0,8,28,1.9,15.8,87.50%,7.4,91,310,3,20,14,3.4,20.7,6.1,119,4.6,547,22.33,119.13,5.33,1.07,6.60,5.33,49.87,9.35,0.27,0.13
DeAndrew White,0,28,9,0,4,2,20,10,0,1,12,0.2,2.2,50.00%,5,,,,0,,,,,2,10,20,1.27,11.87,9.37,0.00,21.53,12.73,157.27,12.35,0.80,0.13
Dede Westbrook,4.1,26,14,10,93,59,588,10,2,26,39,4.2,42,63.40%,6.3,5,27,0,0,8,5.4,1.9,0.4,64,9.6,615,0.67,4.07,6.10,0.07,17.67,10.93,170.00,15.55,1.13,0.07
Deebo Samuel,4.7,23,14,10,76,52,700,13.5,3,28,42,3.7,50,68.40%,9.2,12,126,2,4,31,10.5,9,0.9,64,12.9,826,0.73,2.93,4.00,0.00,17.60,11.93,164.93,13.82,1.00,0.20
Demarcus Robinson,4.1,25,15,10,53,31,425,13.7,3,18,44,2.1,28.3,58.50%,8,,,,0,,,,,31,13.7,425,0.53,5.93,11.12,0.00,17.00,10.53,136.40,12.95,0.87,0.07
Demetrius Harris,2.3,28,14,5,26,15,149,9.9,3,10,23,1.1,10.6,57.70%,5.7,,,,0,,,,,15,9.9,149,0.00,0.00,0.00,0.00,7.80,5.93,72.47,12.21,1.00,0.07
Deon Cain,0,23,12,6,20,9,124,13.8,0,7,35,0.8,10.3,45.00%,6.2,,,,0,,,,,9,13.8,124,0.53,4.33,8.12,0.07,20.60,12.40,136.27,10.99,0.40,0.40
Derek Carrier,1.5,29,15,4,18,12,104,8.7,1,4,25,0.8,6.9,66.70%,5.8,1,27,0,1,27,27,1.8,0.1,13,10.1,131,0.07,0.27,4.00,0.00,6.00,4.20,51.20,12.19,0.47,0.00
Derek Watt,0,27,15,2,5,3,32,10.7,0,1,21,0.2,2.1,60.00%,6.4,7,10,1,6,3,1.4,0.7,0.5,10,4.2,42,22.13,96.27,4.35,0.47,6.53,4.67,36.13,7.74,0.27,0.27
DeVante Parker,23.2,26,15,13,117,64,1065,16.6,9,52,51,4.3,71,54.70%,9.1,,,,0,,,,,64,16.6,1065,0.33,1.73,5.20,0.00,19.60,13.13,186.47,14.20,1.47,0.13
Devin Singletary,8.9,22,12,8,41,29,194,6.7,2,5,49,2.4,16.2,70.70%,4.7,151,775,2,37,38,5.1,64.6,12.6,180,5.4,969,23.40,87.80,3.75,0.27,7.00,4.87,36.67,7.53,0.13,0.27
Devonta Freeman,7.5,27,13,13,67,57,395,6.9,4,16,28,4.4,30.4,85.10%,5.9,166,598,2,27,28,3.6,46,12.8,223,4.5,993,19.27,80.87,4.20,0.40,5.53,3.87,24.67,6.38,0.00,0.33
Devontae Booker,0.5,27,15,0,7,4,40,10,0,1,25,0.3,2.7,57.10%,5.7,2,9,0,0,5,4.5,0.6,0.1,6,8.2,49,22.20,108.87,4.90,0.60,8.00,5.67,55.47,9.79,0.33,0.20
Dion Lewis,9.1,29,15,1,32,25,164,6.6,1,7,24,1.7,10.9,78.10%,5.1,53,202,0,6,17,3.8,13.5,3.5,78,4.7,366,20.67,90.87,4.40,0.40,8.07,6.87,58.93,8.58,0.53,0.07
Diontae Johnson,9.2,23,15,11,85,55,626,11.4,5,29,45,3.7,41.7,64.70%,7.4,4,41,0,2,17,10.3,2.7,0.3,59,11.3,667,0.53,4.33,8.12,0.07,20.60,12.40,136.27,10.99,0.40,0.40
Diontae Spencer,0,27,15,1,8,6,31,5.2,0,1,20,0.4,2.1,75.00%,3.9,2,14,0,0,9,7,0.9,0.1,8,5.6,45,0.40,3.33,8.33,0.00,17.20,9.53,122.40,12.84,0.67,0.07
Dontrell Hilliard,0,24,14,0,15,12,92,7.7,0,4,19,0.9,6.6,80.00%,6.1,13,49,2,3,11,3.8,3.5,0.9,25,5.6,141,23.27,99.73,4.29,0.53,7.20,6.07,50.93,8.40,0.33,0.13
Dontrelle Inman,4.5,30,6,1,18,11,175,15.9,0,9,28,1.8,29.2,61.10%,9.7,,,,0,,,,,11,15.9,175,1.27,13.80,10.89,0.07,21.20,12.67,175.80,13.88,1.20,0.13
Duke Johnson,4.3,26,15,2,56,39,365,9.4,3,15,21,2.6,24.3,69.60%,6.5,79,398,1,16,40,5,26.5,5.3,118,6.5,763,21.60,87.07,4.03,0.80,8.20,6.33,46.87,7.40,0.20,0.13
Durham Smythe,0,24,15,13,11,6,57,9.5,0,2,24,0.4,3.8,54.50%,5.2,,,,0,,,,,6,9.5,57,0.07,0.13,2.00,0.00,6.80,4.40,47.33,10.76,0.47,0.00
Dwayne Washington,2,25,15,0,1,1,6,6,0,0,6,0.1,0.4,100.00%,6,6,58,0,2,31,9.7,3.9,0.4,7,9.1,64,20.13,83.87,4.17,0.27,7.80,6.73,45.33,6.73,0.13,0.27
Elijhaa Penny,-0.2,26,15,1,4,2,9,4.5,0,0,9,0.1,0.6,50.00%,2.3,15,39,0,2,6,2.6,2.6,1,17,2.8,48,27.20,121.07,4.45,0.73,5.40,4.53,39.33,8.68,0.33,0.07
Emmanuel Sanders,2.9,32,16,15,93,63,844,13.4,5,39,75,3.9,52.8,67.70%,9.1,,,,0,,,,,63,13.4,844,0.73,2.93,4.00,0.00,17.60,11.93,164.93,13.82,1.00,0.20
Frank Gore,1.5,36,15,7,12,10,84,8.4,0,4,18,0.7,5.6,83.30%,7,160,573,2,29,41,3.6,38.2,10.7,170,3.9,657,23.40,87.80,3.75,0.27,7.00,4.87,36.67,7.53,0.13,0.27
Fred Brown,0,26,12,1,3,2,21,10.5,0,1,16,0.2,1.8,66.70%,7,,,,0,,,,,2,10.5,21,0.40,3.33,8.33,0.00,17.20,9.53,122.40,12.84,0.67,0.07
Geronimo Allison,3.9,25,15,6,51,31,270,8.7,2,15,31,2.1,18,60.80%,5.3,1,7,0,0,7,7,0.5,0.1,32,8.7,277,0.20,1.13,5.67,0.00,18.93,11.47,147.87,12.90,0.60,0.13
Giovani Bernard,5.7,28,15,2,42,30,234,7.8,0,7,35,2,15.6,71.40%,5.6,50,166,0,10,25,3.3,11.1,3.3,80,5,400,18.93,78.67,4.15,0.07,6.13,4.40,31.33,7.12,0.13,0.27
Golden Tate,12.1,31,10,10,77,44,608,13.8,5,27,64,4.4,60.8,57.10%,7.9,1,16,0,1,16,16,1.6,0.1,45,13.9,624,0.53,1.80,3.38,0.00,20.80,12.33,179.00,14.51,1.80,0.00
Greg Ward,19.1,24,6,2,33,22,211,9.6,1,13,38,3.7,35.2,66.70%,6.4,1,5,0,0,5,5,0.8,0.2,23,9.4,216,0.73,3.93,5.36,0.07,16.87,11.67,142.27,12.19,1.20,0.13
Gus Edwards,3.5,24,15,0,6,6,43,7.2,0,2,10,0.4,2.9,100.00%,7.2,112,581,2,39,63,5.2,38.7,7.5,118,5.3,624,21.27,67.53,3.18,0.67,7.47,5.73,45.33,7.91,0.13,0.07
Hale Hentges,0,23,10,4,7,4,41,10.3,1,3,22,0.4,4.1,57.10%,5.9,,,,0,,,,,4,10.3,41,0.00,0.00,0.00,0.00,5.67,3.80,38.87,10.23,0.27,0.07
Hayden Hurst,2.9,26,15,4,37,28,314,11.2,2,14,61,1.9,20.9,75.70%,8.5,,,,0,,,,,28,11.2,314,0.00,0.27,0.00,0.00,6.20,3.93,41.40,10.53,0.20,0.00
Hunter Henry,2.9,25,11,11,70,50,610,12.2,4,33,30,4.5,55.5,71.40%,8.7,,,,0,,,,,50,12.2,610,0.33,0.33,1.00,0.00,8.47,5.53,51.73,9.35,0.07,0.13
Ian Thomas,4.3,23,15,3,25,15,124,8.3,1,9,19,1,8.3,60.00%,5,,,,0,,,,,15,8.3,124,0.00,0.00,0.00,0.00,8.73,6.00,67.53,11.26,0.40,0.07
Irv Smith Jr.,8.8,21,15,7,45,35,300,8.6,2,16,29,2.3,20,77.80%,6.7,,,,0,,,,,35,8.6,300,0.00,0.00,0.00,0.00,5.93,4.07,44.53,10.95,0.40,0.00
Isaac Nauta,2,22,5,0,3,2,13,6.5,0,1,10,0.4,2.6,66.70%,4.3,,,,0,,,,,2,6.5,13,0.00,0.00,0.00,0.00,7.93,5.00,59.93,11.99,0.47,0.00
Isaiah Ford,5.1,23,7,0,26,16,190,11.9,0,12,28,2.3,27.1,61.50%,7.3,,,,0,,,,,16,11.9,190,0.33,1.73,5.20,0.00,19.60,13.13,186.47,14.20,1.47,0.13
Isaiah McKenzie,0,24,14,7,34,25,247,9.9,1,11,46,1.8,17.6,73.50%,7.3,6,19,0,2,10,3.2,1.4,0.4,31,8.6,266,0.33,2.60,7.80,0.00,18.80,11.07,145.73,13.17,0.87,0.20
J.D. McKissic,2.9,26,15,3,40,33,229,6.9,1,7,26,2.2,15.3,82.50%,5.7,38,205,0,8,44,5.4,13.7,2.5,71,6.1,434,18.13,54.67,3.01,0.53,7.27,5.40,31.00,5.74,0.07,0.40
J.P. Holtz,0.9,26,14,6,8,7,91,13,0,4,30,0.5,6.5,87.50%,11.4,,,,0,,,,,7,13,91,0.00,0.00,0.00,0.00,6.93,4.93,56.33,11.42,0.40,0.13
Jack Doyle,4.1,29,15,15,68,42,442,10.5,4,29,23,2.8,29.5,61.80%,6.5,,,,0,,,,,42,10.5,442,0.07,0.00,0.00,0.00,6.40,4.60,49.87,10.84,0.33,0.07
Jacob Hollister,5.3,26,10,2,51,37,324,8.8,3,15,22,3.7,32.4,72.50%,6.4,,,,0,,,,,37,8.8,324,0.00,0.00,0.00,0.00,5.07,3.40,44.47,13.08,0.20,0.00
Jaeden Graham,0,24,15,0,10,9,149,16.6,1,7,53,0.6,9.9,90.00%,14.9,,,,0,,,,,9,16.6,149,0.00,0.00,0.00,0.00,6.07,4.07,34.80,8.56,0.40,0.07
Jake Kumerow,5.9,27,13,4,19,11,212,19.3,1,8,49,0.8,16.3,57.90%,11.2,,,,0,,,,,11,19.3,212,0.20,1.13,5.67,0.00,18.93,11.47,147.87,12.90,0.60,0.13
Jakobi Meyers,0,23,14,1,41,26,359,13.8,0,17,35,1.9,25.6,63.40%,8.8,,,,0,,,,,26,13.8,359,1.33,7.00,5.25,0.00,17.33,10.47,158.67,15.16,0.73,0.07
Jalen Richard,5.6,26,15,0,41,34,284,8.4,0,14,31,2.3,18.9,82.90%,6.9,36,125,0,10,13,3.5,8.3,2.4,70,5.8,409,22.33,119.13,5.33,1.07,6.60,5.33,49.87,9.35,0.27,0.13
Jamaal Williams,4.3,24,14,2,45,39,253,6.5,5,16,17,2.8,18.1,86.70%,5.6,107,460,1,23,45,4.3,32.9,7.6,146,4.9,713,23.07,84.67,3.67,0.93,7.20,5.47,38.40,7.02,0.13,0.07
James Conner,15.1,24,10,10,38,34,251,7.4,3,14,26,3.4,25.1,89.50%,6.6,116,464,4,26,25,4,46.4,11.6,150,4.8,715,19.93,89.27,4.48,0.60,7.47,5.47,42.33,7.74,0.20,0.13
James Washington,13.3,23,14,9,77,44,735,16.7,3,31,79,3.1,52.5,57.10%,9.5,,,,0,,,,,44,16.7,735,0.53,4.33,8.12,0.07,20.60,12.40,136.27,10.99,0.40,0.40
James White,15.2,27,14,1,92,69,612,8.9,4,29,59,4.9,43.7,75.00%,6.7,65,259,1,15,32,4,18.5,4.6,134,6.5,871,24.87,115.73,4.65,0.80,5.87,4.80,44.20,9.21,0.27,0.20
Jamison Crowder,27,26,15,11,112,70,767,11,5,37,41,4.7,51.1,62.50%,6.8,1,4,0,0,4,4,0.3,0.1,71,10.9,771,0.47,3.73,8.00,0.00,22.60,13.33,166.27,12.47,0.73,0.27
Jared Cook,9.4,32,13,7,63,41,661,16.1,8,30,61,3.2,50.8,65.10%,10.5,,,,0,,,,,41,16.1,661,0.00,0.00,0.00,0.00,7.33,5.33,51.87,9.73,0.40,0.07
Jarius Wright,1.9,30,15,9,53,26,286,11,0,15,33,1.7,19.1,49.10%,5.4,1,-7,0,0,-7,-7,-0.5,0.1,27,10.3,279,1.27,11.87,9.37,0.00,21.53,12.73,157.27,12.35,0.80,0.13
Jaron Brown,1.9,29,13,4,26,16,220,13.8,2,10,48,1.2,16.9,61.50%,8.5,,,,0,,,,,16,13.8,220,0.40,3.40,8.50,0.07,22.20,14.47,180.60,12.48,0.80,0.07
Jason Moore,0,24,9,0,4,2,43,21.5,0,2,32,0.2,4.8,50.00%,10.8,,,,0,,,,,2,21.5,43,0.60,2.00,3.33,0.00,21.27,14.33,171.60,11.97,1.20,0.27
Jason Witten,13.6,37,15,15,79,59,505,8.6,4,25,33,3.9,33.7,74.70%,6.4,,,,0,,,,,59,8.6,505,0.13,0.60,4.50,0.00,6.53,4.33,52.93,12.22,0.33,0.00
Javon Wims,0,25,15,5,32,15,163,10.9,1,7,37,1,10.9,46.90%,5.1,,,,0,,,,,15,10.9,163,0.47,1.40,3.00,0.00,17.67,10.00,159.13,15.91,0.73,0.07
Javorius Allen,8.8,28,9,0,0,0,0,,0,0,0,0,0,0.00%,,9,32,1,2,19,3.6,3.6,1,9,3.6,32,27.20,121.07,4.45,0.73,5.40,4.53,39.33,8.68,0.33,0.07
Jay Ajayi,0,26,3,0,1,0,0,,0,0,0,0,0,0.00%,0,10,30,0,3,11,3,10,3.3,10,3,30,25.80,119.33,4.63,0.67,7.73,6.07,53.13,8.76,0.27,0.20
Jaylen Samuels,1.4,23,13,4,55,46,289,6.3,1,18,27,3.5,22.2,83.60%,5.3,66,175,1,9,13,2.7,13.5,5.1,112,4.1,464,19.93,89.27,4.48,0.60,7.47,5.47,42.33,7.74,0.20,0.13
Jeff Heuerman,0,27,13,10,20,14,114,8.1,1,9,26,1.1,8.8,70.00%,5.7,,,,0,,,,,14,8.1,114,0.00,0.00,0.00,0.00,9.20,6.20,62.13,10.02,0.27,0.00
Jeff Wilson,0,24,10,0,5,3,34,11.3,1,1,25,0.3,3.4,60.00%,6.8,27,105,4,9,25,3.9,10.5,2.7,30,4.6,139,21.60,88.13,4.08,0.53,7.13,5.33,38.40,7.20,0.27,0.20
Jeremy Sprinkle,3.3,25,15,12,34,23,223,9.7,1,12,23,1.5,14.9,67.60%,6.6,,,,0,,,,,23,9.7,223,0.00,0.00,0.00,0.00,5.67,3.80,38.87,10.23,0.27,0.07
Jesper Horsted,0.8,22,5,1,10,8,87,10.9,1,4,20,1.6,17.4,80.00%,8.7,,,,0,,,,,8,10.9,87,0.00,0.00,0.00,0.00,6.93,4.93,56.33,11.42,0.40,0.13
Jesse James,6.1,25,15,10,24,14,137,9.8,0,8,23,0.9,9.1,58.30%,5.7,,,,0,,,,,14,9.8,137,0.00,0.00,0.00,0.00,7.93,5.00,59.93,11.99,0.47,0.00
Jimmy Graham,1,33,15,9,53,34,398,11.7,3,20,48,2.3,26.5,64.20%,7.5,,,,0,,,,,34,11.7,398,0.00,0.00,0.00,0.00,8.53,6.27,57.73,9.21,0.33,0.00
JJ Arcega-Whiteside,0,23,15,5,22,10,169,16.9,1,7,30,0.7,11.3,45.50%,7.7,,,,0,,,,,10,16.9,169,0.73,3.93,5.36,0.07,16.87,11.67,142.27,12.19,1.20,0.13
JJ Nelson,0,27,2,1,5,4,36,9,1,1,29,2,18,80.00%,7.2,,,,0,,,,,4,9,36,0.80,5.27,6.58,0.00,18.60,11.40,160.60,14.09,0.67,0.07
Joe Mixon,18.6,23,15,14,44,34,273,8,3,13,33,2.3,18.2,77.30%,6.2,252,975,3,50,30,3.9,65,16.8,286,4.4,1248,18.93,78.67,4.15,0.07,6.13,4.40,31.33,7.12,0.13,0.27
John Brown,16.9,29,15,15,115,72,1060,14.7,6,53,53,4.8,70.7,62.60%,9.2,2,7,0,0,4,3.5,0.5,0.1,74,14.4,1067,0.33,2.60,7.80,0.00,18.80,11.07,145.73,13.17,0.87,0.20
John Kelly,0,23,3,0,0,0,0,,0,0,0,0,0,0.00%,,3,9,0,0,6,3,3,1,3,3,9,20.40,81.40,3.99,0.73,7.93,6.13,47.00,7.66,0.13,0.13
John Ross,4.4,25,7,7,51,26,464,17.8,3,20,66,3.7,66.3,51.00%,9.1,2,6,0,0,5,3,0.9,0.3,28,16.8,470,0.33,4.80,14.40,0.07,19.87,9.93,117.60,11.84,0.27,0.20
Johnny Holton,1.9,28,15,3,15,3,21,7,0,1,18,0.2,1.4,20.00%,1.4,1,9,0,1,9,9,0.6,0.1,4,7.5,30,0.53,4.33,8.12,0.07,20.60,12.40,136.27,10.99,0.40,0.40
Johnny Mundt,3.5,25,12,2,6,3,24,8,0,1,9,0.3,2,50.00%,4,,,,0,,,,,3,8,24,0.07,0.13,2.00,0.00,8.87,6.47,62.40,9.65,0.40,0.07
Jon Hilliman,0,24,3,1,4,3,1,0.3,0,0,5,1,0.3,75.00%,0.3,30,91,0,6,10,3,30.3,10,33,2.8,92,27.20,121.07,4.45,0.73,5.40,4.53,39.33,8.68,0.33,0.07
Jonathan Williams,0,25,8,1,5,5,59,11.8,0,3,31,0.6,7.4,100.00%,11.8,49,235,1,13,48,4.8,29.4,6.1,54,5.4,294,18.13,67.20,3.71,0.40,7.20,5.73,34.47,6.01,0.27,0.20
Jonnu Smith,16.7,24,15,13,44,35,439,12.5,3,16,57,2.3,29.3,79.50%,10,3,71,0,2,57,23.7,4.7,0.2,38,13.4,510,0.07,3.80,57.00,0.00,7.47,4.87,58.60,12.04,0.33,0.00
Jordan Akins,2.7,27,15,8,48,31,364,11.7,2,18,53,2.1,24.3,64.60%,7.6,,,,0,,,,,31,11.7,364,0.00,0.00,0.00,0.00,7.27,4.93,56.93,11.54,0.60,0.13
Jordan Wilkins,8.7,25,14,1,11,7,43,6.1,0,1,11,0.5,3.1,63.60%,3.9,51,307,2,12,55,6,21.9,3.6,58,6,350,18.13,67.20,3.71,0.40,7.20,5.73,34.47,6.01,0.27,0.20
Josh Adams,0,23,3,0,0,0,0,,0,0,0,0,0,0.00%,,8,12,0,1,10,1.5,4,2.7,8,1.5,12,18.40,80.60,4.38,0.67,5.00,3.93,29.20,7.42,0.07,0.07
Josh Hill,7.5,29,15,10,30,22,191,8.7,3,11,29,1.5,12.7,73.30%,6.4,,,,0,,,,,22,8.7,191,0.00,0.00,0.00,0.00,7.33,5.33,51.87,9.73,0.40,0.07
Josh Jacobs,12.9,21,13,13,27,20,166,8.3,0,8,28,1.5,12.8,74.10%,6.1,242,1150,7,53,51,4.8,88.5,18.6,262,5,1316,22.33,119.13,5.33,1.07,6.60,5.33,49.87,9.35,0.27,0.13
Josh Reynolds,5.6,24,15,2,42,21,326,15.5,1,15,31,1.4,21.7,50.00%,7.8,5,23,0,2,12,4.6,1.5,0.3,26,13.4,349,0.67,3.27,4.90,0.00,17.67,10.87,135.47,12.47,0.80,0.00
Joshua Perkins,0,26,4,0,7,5,37,7.4,0,3,13,1.3,9.3,71.40%,5.3,,,,0,,,,,5,7.4,37,0.13,0.00,0.00,0.00,7.67,5.47,57.27,10.48,0.60,0.00
Julian Edelman,2.9,33,15,13,146,97,1091,11.2,6,53,44,6.5,72.7,66.40%,7.5,8,27,0,2,9,3.4,1.8,0.5,105,10.6,1118,1.33,7.00,5.25,0.00,17.33,10.47,158.67,15.16,0.73,0.07
Justice Hill,1.5,22,15,0,13,7,60,8.6,0,4,14,0.5,4,53.80%,4.6,48,186,1,8,18,3.9,12.4,3.2,55,4.5,246,21.27,67.53,3.18,0.67,7.47,5.73,45.33,7.91,0.13,0.07
Justin Hardy,0,28,15,1,23,16,155,9.7,0,7,23,1.1,10.3,69.60%,6.7,,,,0,,,,,16,9.7,155,1.13,7.53,6.65,0.07,19.27,11.53,129.13,11.20,1.00,0.27
Justin Jackson,3.7,24,6,0,11,9,22,2.4,0,0,9,1.5,3.7,81.80%,2,28,189,0,8,40,6.8,31.5,4.7,37,5.7,211,22.13,96.27,4.35,0.47,6.53,4.67,36.13,7.74,0.27,0.27
Justin Watson,3.7,24,15,1,22,13,132,10.2,2,9,17,0.9,8.8,59.10%,6,,,,0,,,,,13,10.2,132,0.33,1.73,5.20,0.00,22.47,13.73,188.73,13.74,1.20,0.27
Kaden Smith,6.8,22,8,5,31,23,170,7.4,3,7,32,2.9,21.3,74.20%,5.5,,,,0,,,,,23,7.4,170,0.00,0.00,0.00,0.00,7.13,5.00,57.13,11.43,0.33,0.00
Kalif Raymond,1.2,25,8,1,12,9,170,18.9,1,6,52,1.1,21.3,75.00%,14.2,1,-5,0,0,-5,-5,-0.6,0.1,10,16.5,165,0.40,0.07,0.17,0.00,20.67,12.27,166.47,13.57,1.13,0.00
Kareem Hunt,15.6,24,7,2,40,34,253,7.4,1,14,29,4.9,36.1,85.00%,6.3,41,167,2,8,16,4.1,23.9,5.9,75,5.6,420,23.27,99.73,4.29,0.53,7.20,6.07,50.93,8.40,0.33,0.13
Keelan Cole,10.6,26,15,1,31,21,294,14,2,17,55,1.4,19.6,67.70%,9.5,1,6,0,0,6,6,0.4,0.1,22,13.6,300,0.67,4.07,6.10,0.07,17.67,10.93,170.00,15.55,1.13,0.07
Keelan Doss,2.7,23,8,2,14,11,133,12.1,0,6,31,1.4,16.6,78.60%,9.5,,,,0,,,,,11,12.1,133,0.80,5.27,6.58,0.00,18.60,11.40,160.60,14.09,0.67,0.07
Keith Smith,0,27,15,5,3,1,13,13,0,1,13,0.1,0.9,33.30%,4.3,4,9,0,4,3,2.3,0.6,0.3,5,4.4,22,19.27,80.87,4.20,0.40,5.53,3.87,24.67,6.38,0.00,0.33
Kelvin Harmon,4.2,23,15,7,39,27,332,12.3,0,15,30,1.8,22.1,69.20%,8.5,,,,0,,,,,27,12.3,332,0.73,7.67,10.45,0.13,20.40,11.93,176.00,14.75,1.33,0.00
Kendrick Bourne,2.1,24,15,0,44,30,358,11.9,5,23,30,2,23.9,68.20%,8.1,,,,0,,,,,30,11.9,358,0.73,2.93,4.00,0.00,17.60,11.93,164.93,13.82,1.00,0.20
Kenjon Barner,-0.6,29,13,0,8,6,22,3.7,0,1,13,0.5,1.7,75.00%,2.8,4,28,0,1,12,7,2.2,0.3,10,5,50,19.27,80.87,4.20,0.40,5.53,3.87,24.67,6.38,0.00,0.33
Kenny Golladay,7.4,26,15,15,112,62,1118,18,11,49,75,4.1,74.5,55.40%,10,,,,0,,,,,62,18,1118,0.60,4.33,7.22,0.07,24.67,14.73,197.87,13.43,1.40,0.13
Kenny Stills,18.5,27,13,5,55,40,561,14,4,27,45,3.1,43.2,72.70%,10.2,,,,0,,,,,40,14,561,0.60,2.67,4.44,0.00,19.60,12.87,166.93,12.97,0.80,0.07
Kenyan Drake,39.6,25,13,9,64,47,322,6.9,0,14,26,3.6,24.8,73.40%,5,158,757,7,43,80,4.8,58.2,12.2,205,5.3,1079,21.80,106.53,4.89,0.80,5.87,4.67,42.87,9.19,0.27,0.20
Kerrith Whyte,0.5,23,5,0,1,1,9,9,0,1,9,0.2,1.8,100.00%,9,21,121,0,5,21,5.8,24.2,4.2,22,5.9,130,19.93,89.27,4.48,0.60,7.47,5.47,42.33,7.74,0.20,0.13
KhaDarel Hodge,0,24,15,1,8,3,57,19,0,2,41,0.2,3.8,37.50%,7.1,,,,0,,,,,3,19,57,0.33,2.80,8.40,0.00,20.33,13.87,170.33,12.28,0.93,0.07
Khari Blasingame,1,23,5,2,4,3,47,15.7,0,2,24,0.6,9.4,75.00%,11.8,,,,0,,,,,3,15.7,47,20.67,90.87,4.40,0.40,8.07,6.87,58.93,8.58,0.53,0.07
Kyle Rudolph,7.8,30,15,15,48,39,367,9.4,6,24,32,2.6,24.5,81.30%,7.6,,,,0,,,,,39,9.4,367,0.00,0.00,0.00,0.00,5.93,4.07,44.53,10.95,0.40,0.00
Lance Kendricks,0,31,11,1,7,3,50,16.7,0,3,24,0.3,4.5,42.90%,7.1,,,,0,,,,,3,16.7,50,0.33,0.33,1.00,0.00,8.47,5.53,51.73,9.35,0.07,0.13
Laquon Treadwell,0,24,12,0,14,9,184,20.4,1,8,58,0.8,15.3,64.30%,13.1,,,,0,,,,,9,20.4,184,0.53,2.00,3.75,0.00,15.47,11.07,129.33,11.69,0.67,0.00
Larry Fitzgerald,7.2,36,15,15,102,71,759,10.7,4,39,54,4.7,50.6,69.60%,7.4,,,,0,,,,,71,10.7,759,0.87,7.13,8.23,0.00,18.47,11.27,144.00,12.78,0.73,0.07
Latavius Murray,6.9,29,15,7,42,33,221,6.7,1,8,30,2.2,14.7,78.60%,5.3,129,576,5,35,30,4.5,38.4,8.6,162,4.9,797,20.13,83.87,4.17,0.27,7.80,6.73,45.33,6.73,0.13,0.27
Le'Veon Bell,10.8,27,14,14,73,61,425,7,1,19,23,4.4,30.4,83.60%,5.8,229,748,3,31,19,3.3,53.4,16.4,290,4,1173,18.40,80.60,4.38,0.67,5.00,3.93,29.20,7.42,0.07,0.07
Lee Smith,0,32,15,5,5,4,31,7.8,1,2,9,0.3,2.1,80.00%,6.2,,,,0,,,,,4,7.8,31,0.00,0.00,0.00,0.00,5.93,4.13,41.87,10.13,0.53,0.00
Leonard Fournette,12.3,24,15,15,100,76,522,6.9,0,23,27,5.1,34.8,76.00%,5.2,265,1152,3,55,81,4.3,76.8,17.7,341,4.9,1674,20.87,81.53,3.91,0.73,7.40,5.80,51.47,8.87,0.40,0.00
LeSean McCoy,1.6,31,13,9,34,28,181,6.5,1,6,23,2.2,13.9,82.40%,5.3,101,465,4,24,39,4.6,35.8,7.8,129,5,646,23.73,94.00,3.96,0.47,6.53,5.20,34.80,6.69,0.13,0.20
Levine Toilolo,0,28,12,0,2,2,10,5,0,0,8,0.2,0.8,100.00%,5,,,,0,,,,,2,5,10,0.00,0.00,0.00,0.00,7.60,4.87,56.00,11.51,0.33,0.00
Logan Thomas,0,28,15,3,25,15,158,10.5,1,10,17,1,10.5,60.00%,6.3,,,,0,,,,,15,10.5,158,0.00,0.00,0.00,0.00,7.93,5.00,59.93,11.99,0.47,0.00
Luke Stocker,1.9,31,14,9,13,7,43,6.1,0,1,18,0.5,3.1,53.80%,3.3,,,,0,,,,,7,6.1,43,0.00,0.00,0.00,0.00,6.07,4.07,34.80,8.56,0.40,0.07
Mack Hollins,0,26,15,3,23,10,125,12.5,0,7,20,0.7,8.3,43.50%,5.4,,,,0,,,,,10,12.5,125,0.33,1.73,5.20,0.00,19.60,13.13,186.47,14.20,1.47,0.13
Malcolm Brown,0,26,13,1,5,1,10,10,0,0,10,0.1,0.8,20.00%,2,60,229,4,14,17,3.8,17.6,4.6,61,3.9,239,20.40,81.40,3.99,0.73,7.93,6.13,47.00,7.66,0.13,0.13
Malik Turner,5.6,23,15,3,22,15,245,16.3,1,10,33,1,16.3,68.20%,11.1,,,,0,,,,,15,16.3,245,0.40,3.40,8.50,0.07,22.20,14.47,180.60,12.48,0.80,0.07
Marcedes Lewis,1.6,35,15,11,18,14,144,10.3,1,7,25,0.9,9.6,77.80%,8,,,,0,,,,,14,10.3,144,0.00,0.00,0.00,0.00,8.53,6.27,57.73,9.21,0.33,0.00
Marcell Ateman,0,25,10,0,3,2,70,35,0,2,36,0.2,7,66.70%,23.3,,,,0,,,,,2,35,70,0.80,5.27,6.58,0.00,18.60,11.40,160.60,14.09,0.67,0.07
Marcus Johnson,5.7,25,7,5,29,15,246,16.4,2,10,50,2.1,35.1,51.70%,8.5,,,,0,,,,,15,16.4,246,1.27,13.80,10.89,0.07,21.20,12.67,175.80,13.88,1.20,0.13
Marlon Mack,1.9,23,13,11,16,14,82,5.9,0,2,14,1.1,6.3,87.50%,5.1,232,1014,6,62,63,4.4,78,17.8,246,4.5,1096,18.13,67.20,3.71,0.40,7.20,5.73,34.47,6.01,0.27,0.20
Marquez Valdes-Scantling,0,25,15,9,49,24,433,18,2,13,74,1.6,28.9,49.00%,8.8,2,9,0,0,9,4.5,0.6,0.1,26,17,442,0.20,1.13,5.67,0.00,18.93,11.47,147.87,12.90,0.60,0.13
Marquise Brown,14.5,22,13,10,69,44,569,12.9,7,24,83,3.4,43.8,63.80%,8.2,,,,0,,,,,44,12.9,569,0.47,2.20,4.71,0.00,20.87,13.13,164.20,12.50,1.33,0.13
Matt Breida,1.7,24,12,5,21,19,120,6.3,1,6,17,1.6,10,90.50%,5.7,119,607,1,23,83,5.1,50.6,9.9,138,5.3,727,21.60,88.13,4.08,0.53,7.13,5.33,38.40,7.20,0.27,0.20
Matt LaCosse,5.2,27,10,7,19,13,131,10.1,1,6,24,1.3,13.1,68.40%,6.9,,,,0,,,,,13,10.1,131,0.13,0.47,3.50,0.00,6.27,4.40,53.20,12.09,0.40,0.07
Maxx Williams,1.4,25,15,9,17,14,179,12.8,1,10,28,0.9,11.9,82.40%,10.5,,,,0,,,,,14,12.8,179,0.13,1.87,14.00,0.00,6.33,4.20,49.80,11.86,0.60,0.00
Melvin Gordon,7.4,26,11,10,48,36,220,6.1,1,9,25,3.3,20,75.00%,4.6,148,566,7,35,24,3.8,51.5,13.5,184,4.3,786,22.13,96.27,4.35,0.47,6.53,4.67,36.13,7.74,0.27,0.27
Michael Crabtree,0,32,2,1,5,4,22,5.5,0,0,9,2,11,80.00%,4.4,,,,0,,,,,4,5.5,22,0.87,7.13,8.23,0.00,18.47,11.27,144.00,12.78,0.73,0.07
Michael Gallup,1.6,23,13,11,106,61,1009,16.5,3,47,62,4.7,77.6,57.50%,9.5,,,,0,,,,,61,16.5,1009,0.53,1.80,3.38,0.07,19.93,12.53,151.60,12.10,0.80,0.27
Michael Walker,0,23,7,0,3,2,15,7.5,0,1,9,0.3,2.1,66.70%,5,,,,0,,,,,2,7.5,15,0.67,4.07,6.10,0.07,17.67,10.93,170.00,15.55,1.13,0.07
Mike Boone,17.6,24,15,1,1,1,5,5,0,0,5,0.1,0.3,100.00%,5,32,125,2,4,24,3.9,8.3,2.1,33,3.9,130,23.07,94.20,4.08,0.80,7.07,5.60,40.07,7.15,0.27,0.00
Mike Davis,0,26,11,1,8,7,22,3.1,0,1,7,0.6,2,87.50%,2.8,11,25,0,0,8,2.3,2.3,1,18,2.6,47,19.27,82.27,4.27,1.07,6.80,5.53,49.67,8.98,0.07,0.33
Mike Gesicki,8.7,24,15,5,82,47,536,11.4,4,23,34,3.1,35.7,57.30%,6.5,,,,0,,,,,47,11.4,536,0.07,0.13,2.00,0.00,6.80,4.40,47.33,10.76,0.47,0.00
Mike Thomas,1.5,25,15,0,5,2,14,7,0,1,9,0.1,0.9,40.00%,2.8,,,,0,,,,,2,7,14,0.67,3.27,4.90,0.00,17.67,10.87,135.47,12.47,0.80,0.00
Mike Williams,17.1,25,14,14,85,47,963,20.5,2,39,56,3.4,68.8,55.30%,11.3,1,2,0,0,2,2,0.1,0.1,48,20.1,965,0.60,2.00,3.33,0.00,21.27,14.33,171.60,11.97,1.20,0.27
Miles Boykin,7.5,23,15,10,20,13,198,15.2,3,10,50,0.9,13.2,65.00%,9.9,,,,0,,,,,13,15.2,198,0.47,2.20,4.71,0.00,20.87,13.13,164.20,12.50,1.33,0.13
Miles Sanders,35.2,22,15,10,58,47,510,10.9,3,19,45,3.1,34,81.00%,8.8,170,766,3,28,65,4.5,51.1,11.3,217,5.9,1276,25.80,119.33,4.63,0.67,7.73,6.07,53.13,8.76,0.27,0.20
Mo Alie-Cox,0,26,15,2,10,7,78,11.1,0,4,21,0.5,5.2,70.00%,7.8,,,,0,,,,,7,11.1,78,0.07,0.00,0.00,0.00,6.40,4.60,49.87,10.84,0.33,0.07
Mohamed Sanu,3.3,30,14,11,84,56,485,8.7,2,28,28,4,34.6,66.70%,5.8,3,11,0,1,8,3.7,0.8,0.2,59,8.4,496,1.33,7.00,5.25,0.00,17.33,10.47,158.67,15.16,0.73,0.07
MyCole Pruitt,0,27,15,10,6,4,77,19.3,0,2,42,0.3,5.1,66.70%,12.8,,,,0,,,,,4,19.3,77,0.07,3.80,57.00,0.00,7.47,4.87,58.60,12.04,0.33,0.00
Myles Gaskin,9.2,22,7,0,12,7,51,7.3,0,2,20,1,7.3,58.30%,4.3,36,133,1,7,27,3.7,19,5.1,43,4.3,184,24.33,96.80,3.98,0.67,7.07,5.53,45.00,8.13,0.00,0.07
Nick Bellore,0,30,13,1,2,2,23,11.5,1,2,20,0.2,1.8,100.00%,11.5,,,,0,,,,,2,11.5,23,23.40,127.27,5.44,1.67,5.07,3.80,23.47,6.18,0.20,0.07
Nick Boyle,0,26,15,14,41,30,315,10.5,2,13,35,2,21,73.20%,7.7,,,,0,,,,,30,10.5,315,0.00,0.27,0.00,0.00,6.20,3.93,41.40,10.53,0.20,0.00
Nick Vannett,9,26,15,7,22,17,166,9.8,0,5,18,1.1,11.1,77.30%,7.5,,,,0,,,,,17,9.8,166,0.00,0.00,0.00,0.00,5.27,3.80,36.20,9.53,0.33,0.00
Noah Fant,7.6,22,15,11,64,39,558,14.3,3,23,75,2.6,37.2,60.90%,8.7,3,-12,0,0,-2,-4,-0.8,0.2,42,13,546,0.00,0.00,0.00,0.00,9.20,6.20,62.13,10.02,0.27,0.00
Nyheim Hines,3.2,23,15,2,53,41,298,7.3,0,15,21,2.7,19.9,77.40%,5.6,45,165,2,13,18,3.7,11,3,86,5.4,463,18.13,67.20,3.71,0.40,7.20,5.73,34.47,6.01,0.27,0.20
O.J. Howard,8.6,25,13,13,53,34,459,13.5,1,23,33,2.6,35.3,64.20%,8.7,,,,0,,,,,34,13.5,459,0.13,2.00,15.00,0.00,6.47,4.60,51.53,11.20,0.33,0.00
Odell Beckham,14.6,27,15,15,127,71,954,13.4,3,41,89,4.7,63.6,55.90%,7.5,3,10,0,1,11,3.3,0.7,0.2,74,13,964,0.33,2.80,8.40,0.00,20.33,13.87,170.33,12.28,0.93,0.07
Olabisi Johnson,3.5,22,15,5,41,28,260,9.3,3,14,23,1.9,17.3,68.30%,6.3,1,6,0,0,6,6,0.4,0.1,29,9.2,266,0.53,2.00,3.75,0.00,15.47,11.07,129.33,11.69,0.67,0.00
Olamide Zaccheaus,0,22,9,0,3,1,93,93,1,1,93,0.1,10.3,33.30%,31,,,,0,,,,,1,93,93,1.13,7.53,6.65,0.07,19.27,11.53,129.13,11.20,1.00,0.27
Patrick DiMarco,0,30,15,4,7,5,41,8.2,0,1,27,0.3,2.7,71.40%,5.9,3,7,0,0,4,2.3,0.5,0.2,8,6,48,23.40,87.80,3.75,0.27,7.00,4.87,36.67,7.53,0.13,0.27
Patrick Laird,7.4,24,14,3,25,19,156,8.2,0,10,21,1.4,11.1,76.00%,6.2,51,147,1,7,18,2.9,10.5,3.6,70,4.3,303,24.33,96.80,3.98,0.67,7.07,5.53,45.00,8.13,0.00,0.07
Paul Perkins,0,25,4,0,1,1,9,9,0,0,9,0.3,2.3,100.00%,9,12,29,0,3,13,2.4,7.3,3,13,2.9,38,18.13,54.67,3.01,0.53,7.27,5.40,31.00,5.74,0.07,0.40
Peyton Barber,6,25,15,7,20,14,90,6.4,1,3,16,0.9,6,70.00%,4.5,148,460,6,23,17,3.1,30.7,9.9,162,3.4,550,24.33,98.53,4.05,0.87,6.93,5.20,54.40,10.46,0.53,0.33
Pharoh Cooper,2.7,24,12,1,31,24,219,9.1,1,9,28,2,18.3,77.40%,7.1,1,2,0,0,2,2,0.2,0.1,25,8.8,221,0.87,7.13,8.23,0.00,18.47,11.27,144.00,12.78,0.73,0.07
Phillip Dorsett,0,26,13,4,50,28,347,12.4,5,16,58,2.2,26.7,56.00%,6.9,3,21,0,1,9,7,1.6,0.2,31,11.9,368,1.33,7.00,5.25,0.00,17.33,10.47,158.67,15.16,0.73,0.07
Phillip Lindsay,3.2,25,15,15,47,35,196,5.6,0,9,36,2.3,13.1,74.50%,4.2,206,958,7,38,40,4.7,63.9,13.7,241,4.8,1154,22.20,108.87,4.90,0.60,8.00,5.67,55.47,9.79,0.33,0.20
Qadree Ollison,6.1,23,7,0,2,1,7,7,0,1,7,0.1,1,50.00%,3.5,18,41,4,5,6,2.3,5.9,2.6,19,2.5,48,19.27,80.87,4.20,0.40,5.53,3.87,24.67,6.38,0.00,0.33
Raheem Mostert,10.9,27,15,0,20,13,164,12.6,2,6,39,0.9,10.9,65.00%,8.2,127,715,6,27,41,5.6,47.7,8.5,140,6.3,879,21.60,88.13,4.08,0.53,7.13,5.33,38.40,7.20,0.27,0.20
Randall Cobb,0.7,29,14,5,77,50,747,14.9,3,37,59,3.6,53.4,64.90%,9.7,3,11,0,0,7,3.7,0.8,0.2,53,14.3,758,0.53,1.80,3.38,0.07,19.93,12.53,151.60,12.10,0.80,0.27
Rashard Higgins,0,25,10,1,11,4,55,13.8,1,3,35,0.4,5.5,36.40%,5,,,,0,,,,,4,13.8,55,0.33,2.80,8.40,0.00,20.33,13.87,170.33,12.28,0.93,0.07
Reggie Bonnafon,0,23,15,0,7,4,18,4.5,0,0,7,0.3,1.2,57.10%,2.6,14,113,1,2,59,8.1,7.5,0.9,18,7.3,131,19.27,82.27,4.27,1.07,6.80,5.53,49.67,8.98,0.07,0.33
Rex Burkhead,13.9,29,12,1,37,26,273,10.5,0,10,32,2.2,22.8,70.30%,7.4,59,254,3,15,33,4.3,21.2,4.9,85,6.2,527,24.87,115.73,4.65,0.80,5.87,4.80,44.20,9.21,0.27,0.20
Richie James,0,24,15,1,10,6,165,27.5,1,5,57,0.4,11,60.00%,16.5,2,-1,0,0,0,-0.5,-0.1,0.1,8,20.5,164,0.73,2.93,4.00,0.00,17.60,11.93,164.93,13.82,1.00,0.20
Ricky Seals-Jones,15.9,24,13,3,22,14,229,16.4,4,10,59,1.1,17.6,63.60%,10.4,,,,0,,,,,14,16.4,229,0.00,0.00,0.00,0.00,7.80,5.93,72.47,12.21,1.00,0.07
Rico Gafford,0,23,3,1,1,1,49,49,1,1,49,0.3,16.3,100.00%,49,,,,0,,,,,1,49,49,0.80,5.27,6.58,0.00,18.60,11.40,160.60,14.09,0.67,0.07
Riley Ridley,3,23,4,0,3,3,15,5,0,1,13,0.8,3.8,100.00%,5,,,,0,,,,,3,5,15,0.47,1.40,3.00,0.00,17.67,10.00,159.13,15.91,0.73,0.07
Robby Anderson,12.6,26,15,14,89,49,761,15.5,5,34,92,3.3,50.7,55.10%,8.6,1,4,0,0,4,4,0.3,0.1,50,15.3,765,0.47,3.73,8.00,0.00,22.60,13.33,166.27,12.47,0.73,0.27
Robert Davis,0,24,5,2,3,2,17,8.5,0,2,11,0.4,3.4,66.70%,5.7,,,,0,,,,,2,8.5,17,0.73,3.93,5.36,0.07,16.87,11.67,142.27,12.19,1.20,0.13
Robert Foster,0,25,12,1,14,3,64,21.3,0,3,24,0.3,5.3,21.40%,4.6,2,29,0,1,22,14.5,2.4,0.2,5,18.6,93,0.33,2.60,7.80,0.00,18.80,11.07,145.73,13.17,0.87,0.20
Robert Tonyan,1.5,25,10,1,12,8,91,11.4,1,4,28,0.8,9.1,66.70%,7.6,,,,0,,,,,8,11.4,91,0.00,0.00,0.00,0.00,8.53,6.27,57.73,9.21,0.33,0.00
Robert Woods,5.7,27,14,14,127,83,1067,12.9,1,51,48,5.9,76.2,65.40%,8.4,16,106,1,5,20,6.6,7.6,1.1,99,11.8,1173,0.67,3.27,4.90,0.00,17.67,10.87,135.47,12.47,0.80,0.00
Ronald Jones,5.9,22,15,8,38,29,299,10.3,0,12,41,1.9,19.9,76.30%,7.9,161,618,6,30,49,3.8,41.2,10.7,190,4.8,917,24.33,98.53,4.05,0.87,6.93,5.20,54.40,10.46,0.53,0.33
Ross Dwelley,0,24,15,6,22,15,91,6.1,2,8,25,1,6.1,68.20%,4.1,,,,0,,,,,15,6.1,91,0.00,0.00,0.00,0.00,7.60,4.87,56.00,11.51,0.33,0.00
Royce Freeman,6.6,23,15,0,49,42,248,5.9,1,10,19,2.8,16.5,85.70%,5.1,130,500,3,22,26,3.8,33.3,8.7,172,4.3,748,22.20,108.87,4.90,0.60,8.00,5.67,55.47,9.79,0.33,0.20
Russell Gage,8.3,23,15,3,61,42,378,9,1,19,19,2.8,25.2,68.90%,6.2,4,12,0,0,6,3,0.8,0.3,46,8.5,390,1.13,7.53,6.65,0.07,19.27,11.53,129.13,11.20,1.00,0.27
Ryquell Armstead,0.1,23,15,0,15,9,92,10.2,1,5,31,0.6,6.1,60.00%,6.1,25,75,0,2,16,3,5,1.7,34,4.9,167,20.87,81.53,3.91,0.73,7.40,5.80,51.47,8.87,0.40,0.00
Sammy Watkins,9.9,26,13,12,88,51,665,13,3,30,68,3.9,51.2,58.00%,7.6,2,12,0,1,11,6,0.9,0.2,53,12.8,677,0.53,5.93,11.12,0.00,17.00,10.53,136.40,12.95,0.87,0.07
Saquon Barkley,30.3,22,12,12,69,49,413,8.4,2,13,65,4.1,34.4,71.00%,6,200,911,5,43,67,4.6,75.9,16.7,249,5.3,1324,27.20,121.07,4.45,0.73,5.40,4.53,39.33,8.68,0.33,0.07
Scott Miller,13.9,22,10,2,26,13,200,15.4,1,5,48,1.3,20,50.00%,7.7,2,16,0,1,18,8,1.6,0.2,15,14.4,216,0.33,1.73,5.20,0.00,22.47,13.73,188.73,13.74,1.20,0.27
Scott Simonson,1.1,27,5,1,2,2,11,5.5,0,1,10,0.4,2.2,100.00%,5.5,,,,0,,,,,2,5.5,11,0.00,0.00,0.00,0.00,7.13,5.00,57.13,11.43,0.33,0.00
Seth Devalve,4.3,26,11,6,17,11,136,12.4,0,7,20,1,12.4,64.70%,8,,,,0,,,,,11,12.4,136,0.07,-0.33,-5.00,0.00,7.20,4.60,57.07,12.41,0.60,0.00
Seth Roberts,15.6,28,15,0,34,21,271,12.9,2,18,33,1.4,18.1,61.80%,8,,,,0,,,,,21,12.9,271,0.47,2.20,4.71,0.00,20.87,13.13,164.20,12.50,1.33,0.13
Sony Michel,11.3,24,15,13,20,12,94,7.8,0,7,19,0.8,6.3,60.00%,4.7,229,838,6,51,26,3.7,55.9,15.3,241,3.9,932,24.87,115.73,4.65,0.80,5.87,4.80,44.20,9.21,0.27,0.20
Spencer Ware,5.5,28,3,1,7,5,22,4.4,0,1,18,1.7,7.3,71.40%,3.1,17,51,0,3,6,3,17,5.7,22,3.3,73,23.73,94.00,3.96,0.47,6.53,5.20,34.80,6.69,0.13,0.20
Stanley Morgan,0,23,11,0,10,3,18,6,0,0,9,0.3,1.6,30.00%,1.8,,,,0,,,,,3,6,18,0.33,4.80,14.40,0.07,19.87,9.93,117.60,11.84,0.27,0.20
Stefon Diggs,12,26,15,15,94,63,1130,17.9,6,41,66,4.2,75.3,67.00%,12,5,61,0,3,27,12.2,4.1,0.3,68,17.5,1191,0.53,2.00,3.75,0.00,15.47,11.07,129.33,11.69,0.67,0.00
Stephen Carlson,0,23,8,5,7,5,51,10.2,1,2,21,0.6,6.4,71.40%,7.3,,,,0,,,,,5,10.2,51,0.00,0.00,0.00,0.00,7.80,5.93,72.47,12.21,1.00,0.07
Sterling Shepard,20.1,26,9,9,73,52,537,10.3,3,27,36,5.8,59.7,71.20%,7.4,6,72,0,3,23,12,8,0.7,58,10.5,609,0.53,1.80,3.38,0.00,20.80,12.33,179.00,14.51,1.80,0.00
Steven Sims,15.5,22,15,1,48,29,229,7.9,3,15,32,1.9,15.3,60.40%,4.8,8,91,1,2,65,11.4,6.1,0.5,37,8.6,320,0.73,7.67,10.45,0.13,20.40,11.93,176.00,14.75,1.33,0.00
T.J. Jones,0,27,3,0,4,3,38,12.7,1,2,28,1,12.7,75.00%,9.5,,,,0,,,,,3,12.7,38,0.53,1.80,3.38,0.00,20.80,12.33,179.00,14.51,1.80,0.00
T.Y. Hilton,6.5,30,9,9,65,42,429,10.2,5,21,35,4.7,47.7,64.60%,6.6,,,,0,,,,,42,10.2,429,1.27,13.80,10.89,0.07,21.20,12.67,175.80,13.88,1.20,0.13
Tajae Sharpe,4.8,25,14,6,33,24,316,13.2,4,19,47,1.7,22.6,72.70%,9.6,,,,0,,,,,24,13.2,316,0.40,0.07,0.17,0.00,20.67,12.27,166.47,13.57,1.13,0.00
Tanner Hudson,2.4,25,8,1,4,2,26,13,0,1,14,0.3,3.3,50.00%,6.5,,,,0,,,,,2,13,26,0.13,2.00,15.00,0.00,6.47,4.60,51.53,11.20,0.33,0.00
Tarik Cohen,15.5,24,15,10,94,70,412,5.9,3,17,31,4.7,27.5,74.50%,4.4,60,193,0,14,13,3.2,12.9,4,130,4.7,605,22.47,105.87,4.71,0.93,8.07,5.93,42.87,7.22,0.07,0.07
Tavon Austin,13.2,29,13,0,22,12,176,14.7,1,8,59,0.9,13.5,54.50%,8,6,47,1,2,20,7.8,3.6,0.5,18,12.4,223,0.53,1.80,3.38,0.07,19.93,12.53,151.60,12.10,0.80,0.27
Ted Ginn,2.3,34,15,9,54,29,411,14.2,2,19,45,1.9,27.4,53.70%,7.6,3,18,0,2,12,6,1.2,0.2,32,13.4,429,0.67,5.73,8.60,0.13,18.00,12.20,162.33,13.31,1.07,0.00
Terry McLaurin,24,23,14,14,93,58,919,15.8,7,43,75,4.1,65.6,62.40%,9.9,,,,0,,,,,58,15.8,919,0.73,7.67,10.45,0.13,20.40,11.93,176.00,14.75,1.33,0.00
Tevin Coleman,4,26,13,10,28,20,173,8.7,1,9,37,1.5,13.3,71.40%,6.2,132,533,6,26,48,4,41,10.2,152,4.6,706,21.60,88.13,4.08,0.53,7.13,5.33,38.40,7.20,0.27,0.20
Tevin Jones,0,27,5,0,10,4,61,15.3,0,1,28,0.8,12.2,40.00%,6.1,,,,0,,,,,4,15.3,61,0.53,4.33,8.12,0.07,20.60,12.40,136.27,10.99,0.40,0.40
Tim Patrick,5.6,26,7,2,29,15,204,13.6,0,13,38,2.1,29.1,51.70%,7,,,,0,,,,,15,13.6,204,0.40,3.33,8.33,0.00,17.20,9.53,122.40,12.84,0.67,0.07
Todd Gurley,20.8,25,14,14,47,29,186,6.4,2,7,23,2.1,13.3,61.70%,4,203,789,12,49,25,3.9,56.4,14.5,232,4.2,975,20.40,81.40,3.99,0.73,7.93,6.13,47.00,7.66,0.13,0.13
Tony Brooks-James,0,25,3,0,0,0,0,,0,0,0,0,0,0.00%,,8,7,0,0,8,0.9,2.3,2.7,8,0.9,7,19.93,89.27,4.48,0.60,7.47,5.47,42.33,7.74,0.20,0.13
Tony Pollard,22.3,22,14,0,18,14,102,7.3,1,4,21,1,7.3,77.80%,5.7,72,395,2,18,44,5.5,28.2,5.1,86,5.8,497,24.00,99.47,4.14,0.73,6.27,4.33,34.87,8.05,0.27,0.00
Travis Homer,0.7,21,15,0,8,6,26,4.3,0,0,10,0.4,1.7,75.00%,3.3,8,52,0,3,29,6.5,3.5,0.5,14,5.6,78,23.40,127.27,5.44,1.67,5.07,3.80,23.47,6.18,0.20,0.07
Trent Sherfield,0,23,15,1,13,4,80,20,0,4,38,0.3,5.3,30.80%,6.2,,,,0,,,,,4,20,80,0.87,7.13,8.23,0.00,18.47,11.27,144.00,12.78,0.73,0.07
Trevon Wesco,0,24,15,1,2,2,47,23.5,0,2,32,0.1,3.1,100.00%,23.5,1,2,0,1,2,2,0.1,0.1,3,16.3,49,0.07,-0.20,-3.00,0.00,5.27,3.33,37.07,11.12,0.20,0.00
Trevor Davis,0,26,13,4,11,8,111,13.9,0,4,28,0.6,8.5,72.70%,10.1,4,73,1,2,60,18.3,5.6,0.3,12,15.3,184,0.33,1.73,5.20,0.00,19.60,13.13,186.47,14.20,1.47,0.13
Trey Edmunds,0,25,10,0,7,6,48,8,0,2,11,0.6,4.8,85.70%,6.9,22,92,0,2,45,4.2,9.2,2.2,28,5,140,19.93,89.27,4.48,0.60,7.47,5.47,42.33,7.74,0.20,0.13
Troy Fumagalli,1.7,24,10,5,7,5,29,5.8,1,1,9,0.5,2.9,71.40%,4.1,,,,0,,,,,5,5.8,29,0.00,0.00,0.00,0.00,9.20,6.20,62.13,10.02,0.27,0.00
Troymaine Pope,0,26,13,0,3,2,14,7,1,1,13,0.2,1.1,66.70%,4.7,10,20,0,0,8,2,1.5,0.8,12,2.8,34,22.13,96.27,4.35,0.47,6.53,4.67,36.13,7.74,0.27,0.27
Ty Johnson,4,22,15,1,29,24,109,4.5,0,4,13,1.6,7.3,82.80%,3.8,60,208,0,8,17,3.5,13.9,4,84,3.8,317,18.13,54.67,3.01,0.53,7.27,5.40,31.00,5.74,0.07,0.40
Ty Montgomery,2,26,15,2,17,13,90,6.9,0,3,21,0.9,6,76.50%,5.3,32,103,0,2,15,3.2,6.9,2.1,45,4.3,193,18.40,80.60,4.38,0.67,5.00,3.93,29.20,7.42,0.07,0.07
Tyler Boyd,5.6,25,15,14,141,85,987,11.6,5,47,47,5.7,65.8,60.30%,7,4,23,0,1,10,5.8,1.5,0.3,89,11.3,1010,0.33,4.80,14.40,0.07,19.87,9.93,117.60,11.84,0.27,0.20
Tyler Conklin,0,24,14,1,9,7,49,7,0,2,20,0.5,3.5,77.80%,5.4,,,,0,,,,,7,7,49,0.00,0.00,0.00,0.00,5.93,4.07,44.53,10.95,0.40,0.00
Tyler Eifert,7.4,29,15,4,61,41,402,9.8,3,22,27,2.7,26.8,67.20%,6.6,,,,0,,,,,41,9.8,402,0.07,0.27,4.00,0.07,5.80,3.80,42.20,11.11,0.27,0.07
Tyler Higbee,23.1,26,14,14,77,61,650,10.7,2,32,33,4.4,46.4,79.20%,8.4,,,,0,,,,,61,10.7,650,0.07,0.13,2.00,0.00,8.87,6.47,62.40,9.65,0.40,0.07
Tyler Kroft,8.4,27,10,2,10,5,66,13.2,1,5,20,0.5,6.6,50.00%,6.6,,,,0,,,,,5,13.2,66,0.00,0.00,0.00,0.00,5.93,4.13,41.87,10.13,0.53,0.00
Tyler Lockett,26,27,15,15,104,76,1006,13.2,7,49,44,5.1,67.1,73.10%,9.7,4,-5,0,0,3,-1.3,-0.3,0.3,80,12.5,1001,0.40,3.40,8.50,0.07,22.20,14.47,180.60,12.48,0.80,0.07
Tyrell Williams,12.5,27,13,11,64,42,651,15.5,6,33,46,3.2,50.1,65.60%,10.2,,,,0,,,,,42,15.5,651,0.80,5.27,6.58,0.00,18.60,11.40,160.60,14.09,0.67,0.07
Ventell Bryant,0,23,11,0,1,1,15,15,1,1,15,0.1,1.4,100.00%,15,,,,0,,,,,1,15,15,0.53,1.80,3.38,0.07,19.93,12.53,151.60,12.10,0.80,0.27
Virgil Green,0,31,14,4,12,9,78,8.7,1,4,15,0.6,5.6,75.00%,6.5,,,,0,,,,,9,8.7,78,0.33,0.33,1.00,0.00,8.47,5.53,51.73,9.35,0.07,0.13
Vyncint Smith,7,23,12,3,27,14,189,13.5,0,9,37,1.2,15.8,51.90%,7,2,32,1,2,19,16,2.7,0.2,16,13.8,221,0.47,3.73,8.00,0.00,22.60,13.33,166.27,12.47,0.73,0.27
Wendell Smallwood,0,25,14,0,13,9,64,7.1,0,4,18,0.6,4.6,69.20%,4.9,19,76,0,4,17,4,5.4,1.4,28,5,140,18.73,67.80,3.62,0.60,7.47,5.53,40.73,7.36,0.07,0.13
Will Fuller,11.1,25,11,11,71,49,670,13.7,3,26,54,4.5,60.9,69.00%,9.4,,,,0,,,,,49,13.7,670,0.60,2.67,4.44,0.00,19.60,12.87,166.93,12.97,0.80,0.07
Willie Snead,2.5,27,15,10,41,28,317,11.3,5,20,50,1.9,21.1,68.30%,7.7,1,2,0,0,2,2,0.1,0.1,29,11,319,0.47,2.20,4.71,0.00,20.87,13.13,164.20,12.50,1.33,0.13
Zach Line,0.4,29,12,2,10,6,36,6,0,1,12,0.5,3,60.00%,3.6,7,20,0,5,5,2.9,1.7,0.6,13,4.3,56,20.13,83.87,4.17,0.27,7.80,6.73,45.33,6.73,0.13,0.27
Zach Pascal,8.4,25,15,12,69,40,597,14.9,5,28,37,2.7,39.8,58.00%,8.7,1,12,0,1,12,12,0.8,0.1,41,14.9,609,1.27,13.80,10.89,0.07,21.20,12.67,175.80,13.88,1.20,0.13
Zay Jones,1.5,24,14,8,43,25,195,7.8,0,9,23,1.8,13.9,58.10%,4.5,1,3,0,0,3,3,0.2,0.1,26,7.6,198,0.67,3.27,4.90,0.00,17.67,10.87,135.47,12.47,0.80,0.00
